module notgate(
    output y,
    input a
   );
assign y = !a;
endmodule